module main

const (
	lp_nothing_playing = "Nothing is playing"
	lp_filter_media = "Filter the Media"
	lp_videos = "Videos"
	lp_music = "Music"
)
